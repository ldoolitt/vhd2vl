
module Scientific(
input wire clk
);

parameter [31:0] exp1=25e6;
parameter [31:0] exp2=25E6;
parameter exp3=25.0e6;




endmodule
